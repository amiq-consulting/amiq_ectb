/******************************************************************************
 * (C) Copyright 2022 AMIQ All Rights Reserved
 *
 * MODULE:    amiq_ectb_pkg
 * DEVICE:
 * PROJECT:
 * AUTHOR:    andvin
 * DATE:      2022 5:32:36 PM
 *
 * ABSTRACT:  You can customize the file content from Window -> Preferences -> DVT -> Code Templates -> "verilog File"
 *
 *******************************************************************************/

package amiq_ectb_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "amiq_ectb_object.svh"
    `include "amiq_ectb_component.svh"
    `include "amiq_ectb_environment.svh"
    `include "amiq_ectb_sequence.svh"
    `include "amiq_ectb_test.svh"
    
endpackage
